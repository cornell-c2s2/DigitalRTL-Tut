`ifndef PROJECT_REGINC_V
`define PROJECT_REGINC_V

//Registered Incrementer in Verilog


module RegIncVRTL(
input         logic clk,
input  [31:0] logic in,

output [31:0] logic out
);

//Place Implementation here

endmodule;

`endif