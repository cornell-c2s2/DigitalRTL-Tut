`ifndef PROJECT_REGINC_V
`define PROJECT_REGINC_V

//Registered Incrementer in Verilog


module RegIncVRTL(
    input  logic        clk,
    input  logic        reset,
    input  logic [31:0] a,
    output logic [31:0] b
);

/////////////////////////////////
// IMPLEMENT YOUR DESIGN HERE
/////////////////////////////////


endmodule

`endif